module finv_init_m (
    input wire [5:0] m,
    output wire [5:0] m_ );

    function [5:0] f(input [5:0] in);
    begin
        case(in)
            6'b000000: f = 6'b000000;
            6'b000001: f = 6'b111110;
            6'b000010: f = 6'b111100;
            6'b000011: f = 6'b111010;
            6'b000100: f = 6'b111000;
            6'b000101: f = 6'b110110;
            6'b000110: f = 6'b110101;
            6'b000111: f = 6'b110011;
            6'b001000: f = 6'b110001;
            6'b001001: f = 6'b110000;
            6'b001010: f = 6'b101110;
            6'b001011: f = 6'b101101;
            6'b001100: f = 6'b101011;
            6'b001101: f = 6'b101010;
            6'b001110: f = 6'b101001;
            6'b001111: f = 6'b100111;
            6'b010000: f = 6'b100110;
            6'b010001: f = 6'b100101;
            6'b010010: f = 6'b100011;
            6'b010011: f = 6'b100010;
            6'b010100: f = 6'b100001;
            6'b010101: f = 6'b100000;
            6'b010110: f = 6'b011111;
            6'b010111: f = 6'b011110;
            6'b011000: f = 6'b011101;
            6'b011001: f = 6'b011100;
            6'b011010: f = 6'b011011;
            6'b011011: f = 6'b011010;
            6'b011100: f = 6'b011001;
            6'b011101: f = 6'b011000;
            6'b011110: f = 6'b010111;
            6'b011111: f = 6'b010110;
            6'b100000: f = 6'b010101;
            6'b100001: f = 6'b010100;
            6'b100010: f = 6'b010011;
            6'b100011: f = 6'b010010;
            6'b100100: f = 6'b010001;
            6'b100101: f = 6'b010001;
            6'b100110: f = 6'b010000;
            6'b100111: f = 6'b001111;
            6'b101000: f = 6'b001110;
            6'b101001: f = 6'b001110;
            6'b101010: f = 6'b001101;
            6'b101011: f = 6'b001100;
            6'b101100: f = 6'b001011;
            6'b101101: f = 6'b001011;
            6'b101110: f = 6'b001010;
            6'b101111: f = 6'b001001;
            6'b110000: f = 6'b001001;
            6'b110001: f = 6'b001000;
            6'b110010: f = 6'b000111;
            6'b110011: f = 6'b000111;
            6'b110100: f = 6'b000110;
            6'b110101: f = 6'b000110;
            6'b110110: f = 6'b000101;
            6'b110111: f = 6'b000100;
            6'b111000: f = 6'b000100;
            6'b111001: f = 6'b000011;
            6'b111010: f = 6'b000011;
            6'b111011: f = 6'b000010;
            6'b111100: f = 6'b000010;
            6'b111101: f = 6'b000001;
            6'b111110: f = 6'b000001;
            6'b111111: f = 6'b000000;
            default: f = 'x;
        endcase
    end
    endfunction

    assign m_ = f(m);
endmodule

module finv_init (
    input wire [31:0] x,
    output wire [31:0] y,
    input wire ready,
    output wire valid,
    input wire clk,
    input wire rstn );

    assign valid = ready;

    wire s = x[31];
    wire [7:0] e = x[30:23];
    wire [22:0] m = x[22:0];

    wire ys = s;
    wire [7:0] ye = 8'd253 - e + (m[22:17] == '0 ? 8'd1 : 8'd0); // Nobody cares big number!!
    wire [22:0] ym;

    finv_init_m finv_init_m0 (m[22:17], ym[22:17]);

    assign ym[16:0] = '0;

    assign y = e == '0 ? 32'b0 : {ys, ye, ym};

endmodule
