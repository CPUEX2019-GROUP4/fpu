module sqrt_init_m (
    input wire [6:0] m,
    output wire [5:0] m_ );

    function [5:0] f(input [6:0] in);
    begin
        case(in)
            7'b0000000: f = 6'b011010;
            7'b0000001: f = 6'b011011;
            7'b0000010: f = 6'b011011;
            7'b0000011: f = 6'b011100;
            7'b0000100: f = 6'b011101;
            7'b0000101: f = 6'b011101;
            7'b0000110: f = 6'b011110;
            7'b0000111: f = 6'b011111;
            7'b0001000: f = 6'b100000;
            7'b0001001: f = 6'b100000;
            7'b0001010: f = 6'b100001;
            7'b0001011: f = 6'b100001;
            7'b0001100: f = 6'b100010;
            7'b0001101: f = 6'b100011;
            7'b0001110: f = 6'b100011;
            7'b0001111: f = 6'b100100;
            7'b0010000: f = 6'b100101;
            7'b0010001: f = 6'b100101;
            7'b0010010: f = 6'b100110;
            7'b0010011: f = 6'b100111;
            7'b0010100: f = 6'b100111;
            7'b0010101: f = 6'b101000;
            7'b0010110: f = 6'b101000;
            7'b0010111: f = 6'b101001;
            7'b0011000: f = 6'b101010;
            7'b0011001: f = 6'b101010;
            7'b0011010: f = 6'b101011;
            7'b0011011: f = 6'b101011;
            7'b0011100: f = 6'b101100;
            7'b0011101: f = 6'b101101;
            7'b0011110: f = 6'b101101;
            7'b0011111: f = 6'b101110;
            7'b0100000: f = 6'b101110;
            7'b0100001: f = 6'b101111;
            7'b0100010: f = 6'b110000;
            7'b0100011: f = 6'b110000;
            7'b0100100: f = 6'b110001;
            7'b0100101: f = 6'b110001;
            7'b0100110: f = 6'b110010;
            7'b0100111: f = 6'b110010;
            7'b0101000: f = 6'b110011;
            7'b0101001: f = 6'b110011;
            7'b0101010: f = 6'b110100;
            7'b0101011: f = 6'b110101;
            7'b0101100: f = 6'b110101;
            7'b0101101: f = 6'b110110;
            7'b0101110: f = 6'b110110;
            7'b0101111: f = 6'b110111;
            7'b0110000: f = 6'b110111;
            7'b0110001: f = 6'b111000;
            7'b0110010: f = 6'b111000;
            7'b0110011: f = 6'b111001;
            7'b0110100: f = 6'b111001;
            7'b0110101: f = 6'b111010;
            7'b0110110: f = 6'b111010;
            7'b0110111: f = 6'b111011;
            7'b0111000: f = 6'b111011;
            7'b0111001: f = 6'b111100;
            7'b0111010: f = 6'b111100;
            7'b0111011: f = 6'b111101;
            7'b0111100: f = 6'b111101;
            7'b0111101: f = 6'b111110;
            7'b0111110: f = 6'b111110;
            7'b0111111: f = 6'b111111;
            7'b1000000: f = 6'b000000;
            7'b1000001: f = 6'b000000;
            7'b1000010: f = 6'b000000;
            7'b1000011: f = 6'b000001;
            7'b1000100: f = 6'b000001;
            7'b1000101: f = 6'b000010;
            7'b1000110: f = 6'b000010;
            7'b1000111: f = 6'b000011;
            7'b1001000: f = 6'b000011;
            7'b1001001: f = 6'b000100;
            7'b1001010: f = 6'b000100;
            7'b1001011: f = 6'b000101;
            7'b1001100: f = 6'b000101;
            7'b1001101: f = 6'b000110;
            7'b1001110: f = 6'b000110;
            7'b1001111: f = 6'b000111;
            7'b1010000: f = 6'b000111;
            7'b1010001: f = 6'b001000;
            7'b1010010: f = 6'b001000;
            7'b1010011: f = 6'b001000;
            7'b1010100: f = 6'b001001;
            7'b1010101: f = 6'b001001;
            7'b1010110: f = 6'b001010;
            7'b1010111: f = 6'b001010;
            7'b1011000: f = 6'b001011;
            7'b1011001: f = 6'b001011;
            7'b1011010: f = 6'b001011;
            7'b1011011: f = 6'b001100;
            7'b1011100: f = 6'b001100;
            7'b1011101: f = 6'b001101;
            7'b1011110: f = 6'b001101;
            7'b1011111: f = 6'b001101;
            7'b1100000: f = 6'b001110;
            7'b1100001: f = 6'b001110;
            7'b1100010: f = 6'b001111;
            7'b1100011: f = 6'b001111;
            7'b1100100: f = 6'b010000;
            7'b1100101: f = 6'b010000;
            7'b1100110: f = 6'b010000;
            7'b1100111: f = 6'b010001;
            7'b1101000: f = 6'b010001;
            7'b1101001: f = 6'b010001;
            7'b1101010: f = 6'b010010;
            7'b1101011: f = 6'b010010;
            7'b1101100: f = 6'b010011;
            7'b1101101: f = 6'b010011;
            7'b1101110: f = 6'b010011;
            7'b1101111: f = 6'b010100;
            7'b1110000: f = 6'b010100;
            7'b1110001: f = 6'b010101;
            7'b1110010: f = 6'b010101;
            7'b1110011: f = 6'b010101;
            7'b1110100: f = 6'b010110;
            7'b1110101: f = 6'b010110;
            7'b1110110: f = 6'b010110;
            7'b1110111: f = 6'b010111;
            7'b1111000: f = 6'b010111;
            7'b1111001: f = 6'b011000;
            7'b1111010: f = 6'b011000;
            7'b1111011: f = 6'b011000;
            7'b1111100: f = 6'b011001;
            7'b1111101: f = 6'b011001;
            7'b1111110: f = 6'b011001;
            7'b1111111: f = 6'b011010;
            default: f = 'x;
        endcase
    end
    endfunction

    assign m_ = f(m);
endmodule

module sqrt_init (
    input wire [31:0] x,
    output wire [31:0] y,
    input wire ready,
    output wire valid,
    input wire clk,
    input wire rstn );

    assign valid = ready;

    wire s = x[31];
    wire [7:0] e = x[30:23];
    wire [22:0] m = x[22:0];

    wire ys = s;
    wire [7:0] ye = ((e - 8'd1) >> 1) + 8'd64;
    wire [22:0] ym;

    sqrt_init_m sqrt_init_m0({e[0], m[22:17]}, ym[22:17]);

    assign ym[16:0] = '0;

    assign y = e == '0 ? 32'b0 : {ys, ye, ym};

endmodule
