module fclt (
    input wire [31:0] x1,
    input wire [31:0] x2,
    output wire y,
    input wire ready,
    output wire valid,
    input wire clk,
    input wire rstn );

    assign valid = ready;

    wire s1 = x1[31];
    wire s2 = x2[31];
    wire [30:0] em1 = x1[30:0];
    wire [30:0] em2 = x2[30:0];

    assign y = (s1 && ~s2) || (s1 && s2 && em1 <= em2) || (~s1 && ~s2 && em1 >= em2);

endmodule
